/*
module int_display(I, );

input I;

always @(*)
    begin
        if(sel == 'h0)
            out = a;
        else if(sel == 'h1)
            out = b;
        else if(sel == 'h2)
            out = c;
        else if(sel == 'h3)
            out = d;
    end*/